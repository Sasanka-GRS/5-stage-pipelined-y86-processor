`timescale 1ns / 1ps
module XOR(a,b,y);
input [63:0] a;
input [63:0] b;
output [63:0] y;

xor(y[0],a[0],b[0]);
xor(y[1],a[1],b[1]);
xor(y[2],a[2],b[2]);
xor(y[3],a[3],b[3]);
xor(y[4],a[4],b[4]);
xor(y[5],a[5],b[5]);
xor(y[6],a[6],b[6]);
xor(y[7],a[7],b[7]);
xor(y[8],a[8],b[8]);
xor(y[9],a[9],b[9]);
xor(y[10],a[10],b[10]);
xor(y[11],a[11],b[11]);
xor(y[12],a[12],b[12]);
xor(y[13],a[13],b[13]);
xor(y[14],a[14],b[14]);
xor(y[15],a[15],b[15]);
xor(y[16],a[16],b[16]);
xor(y[17],a[17],b[17]);
xor(y[18],a[18],b[18]);
xor(y[19],a[19],b[19]);
xor(y[20],a[20],b[20]);
xor(y[21],a[21],b[21]);
xor(y[22],a[22],b[22]);
xor(y[23],a[23],b[23]);
xor(y[24],a[24],b[24]);
xor(y[25],a[25],b[25]);
xor(y[26],a[26],b[26]);
xor(y[27],a[27],b[27]);
xor(y[28],a[28],b[28]);
xor(y[29],a[29],b[29]);
xor(y[30],a[30],b[30]);
xor(y[31],a[31],b[31]);
xor(y[32],a[32],b[32]);
xor(y[33],a[33],b[33]);
xor(y[34],a[34],b[34]);
xor(y[35],a[35],b[35]);
xor(y[36],a[36],b[36]);
xor(y[37],a[37],b[37]);
xor(y[38],a[38],b[38]);
xor(y[39],a[39],b[39]);
xor(y[40],a[40],b[40]);
xor(y[41],a[41],b[41]);
xor(y[42],a[42],b[42]);
xor(y[43],a[43],b[43]);
xor(y[44],a[44],b[44]);
xor(y[45],a[45],b[45]);
xor(y[46],a[46],b[46]);
xor(y[47],a[47],b[47]);
xor(y[48],a[48],b[48]);
xor(y[49],a[49],b[49]);
xor(y[50],a[50],b[50]);
xor(y[51],a[51],b[51]);
xor(y[52],a[52],b[52]);
xor(y[53],a[53],b[53]);
xor(y[54],a[54],b[54]);
xor(y[55],a[55],b[55]);
xor(y[56],a[56],b[56]);
xor(y[57],a[57],b[57]);
xor(y[58],a[58],b[58]);
xor(y[59],a[59],b[59]);
xor(y[60],a[60],b[60]);
xor(y[61],a[61],b[61]);
xor(y[62],a[62],b[62]);
xor(y[63],a[63],b[63]);

endmodule